always@(posedge clk or negedge rst) begin

end
